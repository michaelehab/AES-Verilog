module AES(x,y);
input [128:0] x;
output [128:0] y;
mixColumns(x,y);
//To be edited later. This part was added only as it displayed errors when this top module was empty
endmodule