module AES_Encrypt;
endmodule