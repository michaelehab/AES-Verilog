module sbox;
endmodule