module keyExpansion;
endmodule