module keyExpansion;