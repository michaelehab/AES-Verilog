module inverseShiftRows_tb;

reg [127:0] in;
wire [127:0] out;	


inverseShiftRows m (in,out);


initial begin
	$monitor("input= %H , output= %h",in,out);
	in = 128'h_7ad5fda789ef4e272bca100b3d9ff59f;
end
endmodule