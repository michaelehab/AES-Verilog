module addRoundKey;
endmodule