module subBytes;

endmodule