module AES_Decrypt;
endmodule