module mixColumns();

