module AES;

endmodule