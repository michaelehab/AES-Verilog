module AES_Decrypt;