module shiftRows();
endmodule