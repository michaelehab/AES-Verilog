module shiftRows;
endmodule