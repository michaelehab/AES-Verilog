module sbox;