module shiftRows;