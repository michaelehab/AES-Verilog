module rcon;
endmodule